package wishbone_package;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    //`include "wishbone_interface.sv"
    `include "wishbone_sequence.sv"
    `include "wishbone_sequencer.sv"
    `include "wishbone_driver.sv"
    `include "wishbone_monitor.sv"
    `include "wishbone_agent.sv"
    `include "wishbone_scoreboarder.sv"
    `include "wishbone_env.sv"
    `include "wishbone_test.sv"
endpackage



